(* src = "design.sv:2" *)
module Ram_128B(Address, Data, CS, WE, OE);
  (* src = "design.sv:2" *)
  wire [15:0] _000_;
  (* src = "design.sv:16" *)
  wire [15:0] _001_;
  (* src = "design.sv:16" *)
  wire [15:0] _002_;
  (* src = "design.sv:16" *)
  wire [15:0] _003_;
  (* src = "design.sv:16" *)
  wire [15:0] _004_;
  (* src = "design.sv:16" *)
  wire [15:0] _005_;
  (* src = "design.sv:16" *)
  wire [15:0] _006_;
  (* src = "design.sv:16" *)
  wire [15:0] _007_;
  (* src = "design.sv:16" *)
  wire [15:0] _008_;
  (* src = "design.sv:16" *)
  wire [15:0] _009_;
  (* src = "design.sv:16" *)
  wire [15:0] _010_;
  (* src = "design.sv:16" *)
  wire [15:0] _011_;
  (* src = "design.sv:16" *)
  wire [15:0] _012_;
  (* src = "design.sv:16" *)
  wire [15:0] _013_;
  (* src = "design.sv:16" *)
  wire [15:0] _014_;
  (* src = "design.sv:16" *)
  wire [15:0] _015_;
  (* src = "design.sv:16" *)
  wire [15:0] _016_;
  (* src = "design.sv:16" *)
  wire [15:0] _017_;
  (* src = "design.sv:16" *)
  wire [15:0] _018_;
  (* src = "design.sv:16" *)
  wire [15:0] _019_;
  (* src = "design.sv:16" *)
  wire [15:0] _020_;
  (* src = "design.sv:16" *)
  wire [15:0] _021_;
  (* src = "design.sv:16" *)
  wire [15:0] _022_;
  (* src = "design.sv:16" *)
  wire [15:0] _023_;
  (* src = "design.sv:16" *)
  wire [15:0] _024_;
  (* src = "design.sv:16" *)
  wire [15:0] _025_;
  (* src = "design.sv:16" *)
  wire [15:0] _026_;
  (* src = "design.sv:16" *)
  wire [15:0] _027_;
  (* src = "design.sv:16" *)
  wire [15:0] _028_;
  (* src = "design.sv:16" *)
  wire [15:0] _029_;
  (* src = "design.sv:16" *)
  wire [15:0] _030_;
  (* src = "design.sv:16" *)
  wire [15:0] _031_;
  (* src = "design.sv:16" *)
  wire [15:0] _032_;
  (* src = "design.sv:16" *)
  wire [15:0] _033_;
  (* src = "design.sv:16" *)
  wire [15:0] _034_;
  (* src = "design.sv:16" *)
  wire [15:0] _035_;
  (* src = "design.sv:16" *)
  wire [15:0] _036_;
  (* src = "design.sv:16" *)
  wire [15:0] _037_;
  (* src = "design.sv:16" *)
  wire [15:0] _038_;
  (* src = "design.sv:16" *)
  wire [15:0] _039_;
  (* src = "design.sv:16" *)
  wire [15:0] _040_;
  (* src = "design.sv:16" *)
  wire [15:0] _041_;
  (* src = "design.sv:16" *)
  wire [15:0] _042_;
  (* src = "design.sv:16" *)
  wire [15:0] _043_;
  (* src = "design.sv:16" *)
  wire [15:0] _044_;
  (* src = "design.sv:16" *)
  wire [15:0] _045_;
  (* src = "design.sv:16" *)
  wire [15:0] _046_;
  (* src = "design.sv:16" *)
  wire [15:0] _047_;
  (* src = "design.sv:16" *)
  wire [15:0] _048_;
  (* src = "design.sv:16" *)
  wire [15:0] _049_;
  (* src = "design.sv:16" *)
  wire [15:0] _050_;
  (* src = "design.sv:16" *)
  wire [15:0] _051_;
  (* src = "design.sv:16" *)
  wire [15:0] _052_;
  (* src = "design.sv:16" *)
  wire [15:0] _053_;
  (* src = "design.sv:16" *)
  wire [15:0] _054_;
  (* src = "design.sv:16" *)
  wire [15:0] _055_;
  (* src = "design.sv:16" *)
  wire [15:0] _056_;
  (* src = "design.sv:16" *)
  wire [15:0] _057_;
  (* src = "design.sv:16" *)
  wire [15:0] _058_;
  (* src = "design.sv:16" *)
  wire [15:0] _059_;
  (* src = "design.sv:16" *)
  wire [15:0] _060_;
  (* src = "design.sv:16" *)
  wire [15:0] _061_;
  (* src = "design.sv:16" *)
  wire [15:0] _062_;
  (* src = "design.sv:16" *)
  wire [15:0] _063_;
  (* src = "design.sv:16" *)
  wire [15:0] _064_;
  (* src = "design.sv:16" *)
  wire _065_;
  (* src = "design.sv:16" *)
  wire _066_;
  (* src = "design.sv:16" *)
  wire [15:0] _067_;
  (* src = "design.sv:16" *)
  wire _068_;
  (* src = "design.sv:16" *)
  wire [15:0] _069_;
  (* src = "design.sv:16" *)
  wire [15:0] _070_;
  (* src = "design.sv:16" *)
  wire [15:0] _071_;
  (* src = "design.sv:16" *)
  wire [15:0] _072_;
  (* src = "design.sv:16" *)
  wire [15:0] _073_;
  (* src = "design.sv:16" *)
  wire [15:0] _074_;
  (* src = "design.sv:16" *)
  wire [15:0] _075_;
  (* src = "design.sv:16" *)
  wire [15:0] _076_;
  (* src = "design.sv:16" *)
  wire [15:0] _077_;
  (* src = "design.sv:16" *)
  wire [15:0] _078_;
  (* src = "design.sv:16" *)
  wire [15:0] _079_;
  (* src = "design.sv:16" *)
  wire [15:0] _080_;
  (* src = "design.sv:16" *)
  wire [15:0] _081_;
  (* src = "design.sv:16" *)
  wire [15:0] _082_;
  (* src = "design.sv:16" *)
  wire [15:0] _083_;
  (* src = "design.sv:16" *)
  wire [15:0] _084_;
  (* src = "design.sv:16" *)
  wire [15:0] _085_;
  (* src = "design.sv:16" *)
  wire [15:0] _086_;
  (* src = "design.sv:16" *)
  wire [15:0] _087_;
  (* src = "design.sv:16" *)
  wire [15:0] _088_;
  (* src = "design.sv:16" *)
  wire [15:0] _089_;
  (* src = "design.sv:16" *)
  wire [15:0] _090_;
  (* src = "design.sv:16" *)
  wire [15:0] _091_;
  (* src = "design.sv:16" *)
  wire [15:0] _092_;
  (* src = "design.sv:16" *)
  wire [15:0] _093_;
  (* src = "design.sv:16" *)
  wire [15:0] _094_;
  (* src = "design.sv:16" *)
  wire [15:0] _095_;
  (* src = "design.sv:16" *)
  wire [15:0] _096_;
  (* src = "design.sv:16" *)
  wire [15:0] _097_;
  (* src = "design.sv:16" *)
  wire [15:0] _098_;
  (* src = "design.sv:16" *)
  wire [15:0] _099_;
  (* src = "design.sv:16" *)
  wire [15:0] _100_;
  (* src = "design.sv:16" *)
  wire [15:0] _101_;
  (* src = "design.sv:16" *)
  wire [15:0] _102_;
  (* src = "design.sv:16" *)
  wire [15:0] _103_;
  (* src = "design.sv:16" *)
  wire [15:0] _104_;
  (* src = "design.sv:16" *)
  wire [15:0] _105_;
  (* src = "design.sv:16" *)
  wire [15:0] _106_;
  (* src = "design.sv:16" *)
  wire [15:0] _107_;
  (* src = "design.sv:16" *)
  wire [15:0] _108_;
  (* src = "design.sv:16" *)
  wire [15:0] _109_;
  (* src = "design.sv:16" *)
  wire [15:0] _110_;
  (* src = "design.sv:16" *)
  wire [15:0] _111_;
  (* src = "design.sv:16" *)
  wire [15:0] _112_;
  (* src = "design.sv:16" *)
  wire [15:0] _113_;
  (* src = "design.sv:16" *)
  wire [15:0] _114_;
  (* src = "design.sv:16" *)
  wire [15:0] _115_;
  (* src = "design.sv:16" *)
  wire [15:0] _116_;
  (* src = "design.sv:16" *)
  wire [15:0] _117_;
  (* src = "design.sv:16" *)
  wire [15:0] _118_;
  (* src = "design.sv:16" *)
  wire [15:0] _119_;
  (* src = "design.sv:16" *)
  wire [15:0] _120_;
  (* src = "design.sv:16" *)
  wire [15:0] _121_;
  (* src = "design.sv:16" *)
  wire [15:0] _122_;
  (* src = "design.sv:16" *)
  wire [15:0] _123_;
  (* src = "design.sv:16" *)
  wire [15:0] _124_;
  (* src = "design.sv:16" *)
  wire [15:0] _125_;
  (* src = "design.sv:16" *)
  wire [15:0] _126_;
  (* src = "design.sv:16" *)
  wire [15:0] _127_;
  (* src = "design.sv:16" *)
  wire [15:0] _128_;
  (* src = "design.sv:16" *)
  wire [15:0] _129_;
  (* src = "design.sv:16" *)
  wire [15:0] _130_;
  (* src = "design.sv:16" *)
  wire [15:0] _131_;
  (* src = "design.sv:16" *)
  wire [15:0] _132_;
  (* src = "design.sv:16" *)
  wire [15:0] _133_;
  (* src = "design.sv:17" *)
  wire _134_;
  (* src = "design.sv:21" *)
  wire _135_;
  (* src = "design.sv:30" *)
  wire _136_;
  (* src = "design.sv:14" *)
  wire _137_;
  (* src = "design.sv:17" *)
  wire _138_;
  (* src = "design.sv:21" *)
  wire _139_;
  (* src = "design.sv:21" *)
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire _200_;
  wire _201_;
  wire _202_;
  wire _203_;
  (* src = "design.sv:7" *)
  input [5:0] Address;
  (* src = "design.sv:9" *)
  input CS;
  (* src = "design.sv:8" *)
  inout [15:0] Data;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[0] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[10] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[11] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[12] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[13] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[14] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[15] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[16] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[17] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[18] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[19] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[1] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[20] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[21] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[22] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[23] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[24] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[25] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[26] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[27] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[28] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[29] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[2] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[30] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[31] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[32] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[33] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[34] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[35] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[36] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[37] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[38] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[39] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[3] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[40] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[41] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[42] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[43] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[44] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[45] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[46] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[47] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[48] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[49] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[4] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[50] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[51] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[52] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[53] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[54] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[55] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[56] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[57] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[58] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[59] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[5] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[60] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[61] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[62] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[63] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[6] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[7] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[8] ;
  (* src = "design.sv:2" *)
  wire [15:0] \Mem[9] ;
  (* src = "design.sv:9" *)
  input OE;
  (* src = "design.sv:9" *)
  input WE;
  (* src = "design.sv:12" *)
  wire bug_a;
  assign _134_ = _138_ && (* src = "design.sv:17" *) OE;
  assign _135_ = _139_ && (* src = "design.sv:21" *) _140_;
  assign _136_ = _138_ && (* src = "design.sv:30" *) _137_;
  assign _137_ = ! (* src = "design.sv:14" *) OE;
  assign _138_ = ! (* src = "design.sv:17" *) WE;
  assign _139_ = 1023 < (* src = "design.sv:21" *) Data;
  assign _140_ = Data < (* src = "design.sv:21" *) 2048;
  assign _141_ = Address == 6'b010001;
  assign _142_ = Address == 6'b010000;
  assign _143_ = Address == 6'b001111;
  assign _144_ = Address == 6'b001110;
  assign _145_ = Address == 6'b001101;
  assign _146_ = Address == 6'b001100;
  assign _147_ = Address == 6'b001011;
  assign _148_ = Address == 6'b001010;
  assign _149_ = Address == 6'b001001;
  assign _150_ = Address == 6'b001000;
  assign _151_ = Address == 6'b000111;
  assign _152_ = Address == 6'b000110;
  assign _153_ = Address == 6'b000101;
  assign _154_ = Address == 6'b000100;
  assign _155_ = Address == 6'b000011;
  assign _156_ = Address == 6'b000010;
  assign _157_ = Address == 6'b000001;
  assign _158_ = Address == 6'b000000;
  assign _159_ = Address == 6'b100100;
  assign _160_ = Address == 6'b100011;
  assign _161_ = Address == 6'b100010;
  assign _162_ = Address == 6'b100001;
  assign _163_ = Address == 6'b100000;
  assign _164_ = Address == 6'b011111;
  assign _165_ = Address == 6'b011110;
  assign _166_ = Address == 6'b011101;
  assign _167_ = Address == 6'b011100;
  assign _168_ = Address == 6'b011011;
  assign _169_ = Address == 6'b011010;
  assign _170_ = Address == 6'b011001;
  assign _171_ = Address == 6'b011000;
  assign _172_ = Address == 6'b010111;
  assign _173_ = Address == 6'b010110;
  assign _174_ = Address == 6'b010101;
  assign _175_ = Address == 6'b010100;
  assign _176_ = Address == 6'b010011;
  assign _177_ = Address == 6'b010010;
  assign _178_ = Address == 6'b100101;
  assign _179_ = Address == 6'b100110;
  assign _180_ = Address == 6'b100111;
  assign _181_ = Address == 6'b101000;
  assign _182_ = Address == 6'b101001;
  assign _183_ = Address == 6'b101010;
  assign _184_ = Address == 6'b101011;
  assign _185_ = Address == 6'b101100;
  assign _186_ = Address == 6'b101101;
  assign _187_ = Address == 6'b101110;
  assign _188_ = Address == 6'b101111;
  assign _189_ = Address == 6'b110000;
  assign _190_ = Address == 6'b110001;
  assign _191_ = Address == 6'b110010;
  assign _192_ = Address == 6'b110011;
  assign _193_ = Address == 6'b110100;
  assign _194_ = Address == 6'b110101;
  assign _195_ = Address == 6'b110110;
  assign _196_ = Address == 6'b110111;
  assign _197_ = Address == 6'b111000;
  assign _198_ = Address == 6'b111001;
  assign _199_ = Address == 6'b111010;
  assign _200_ = Address == 6'b111011;
  assign _201_ = Address == 6'b111100;
  assign _202_ = Address == 6'b111101;
  assign _203_ = Address == 6'b111110;
  reg [15:0] _274_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _274_ = _070_;
      default:
        _274_ = _001_;
    endcase
  assign \Mem[0]  = _274_;
  reg [15:0] _275_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _275_ = _071_;
      default:
        _275_ = _002_;
    endcase
  assign \Mem[10]  = _275_;
  reg [15:0] _276_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _276_ = _072_;
      default:
        _276_ = _003_;
    endcase
  assign \Mem[11]  = _276_;
  reg [15:0] _277_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _277_ = _073_;
      default:
        _277_ = _004_;
    endcase
  assign \Mem[12]  = _277_;
  reg [15:0] _278_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _278_ = _074_;
      default:
        _278_ = _005_;
    endcase
  assign \Mem[13]  = _278_;
  reg [15:0] _279_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _279_ = _075_;
      default:
        _279_ = _006_;
    endcase
  assign \Mem[14]  = _279_;
  reg [15:0] _280_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _280_ = _076_;
      default:
        _280_ = _007_;
    endcase
  assign \Mem[15]  = _280_;
  reg [15:0] _281_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _281_ = _077_;
      default:
        _281_ = _008_;
    endcase
  assign \Mem[16]  = _281_;
  reg [15:0] _282_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _282_ = _078_;
      default:
        _282_ = _009_;
    endcase
  assign \Mem[17]  = _282_;
  reg [15:0] _283_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _283_ = _079_;
      default:
        _283_ = _010_;
    endcase
  assign \Mem[18]  = _283_;
  reg [15:0] _284_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _284_ = _080_;
      default:
        _284_ = _011_;
    endcase
  assign \Mem[19]  = _284_;
  reg [15:0] _285_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _285_ = _081_;
      default:
        _285_ = _012_;
    endcase
  assign \Mem[1]  = _285_;
  reg [15:0] _286_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _286_ = _082_;
      default:
        _286_ = _013_;
    endcase
  assign \Mem[20]  = _286_;
  reg [15:0] _287_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _287_ = _083_;
      default:
        _287_ = _014_;
    endcase
  assign \Mem[21]  = _287_;
  reg [15:0] _288_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _288_ = _084_;
      default:
        _288_ = _015_;
    endcase
  assign \Mem[22]  = _288_;
  reg [15:0] _289_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _289_ = _085_;
      default:
        _289_ = _016_;
    endcase
  assign \Mem[23]  = _289_;
  reg [15:0] _290_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _290_ = _086_;
      default:
        _290_ = _017_;
    endcase
  assign \Mem[24]  = _290_;
  reg [15:0] _291_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _291_ = _087_;
      default:
        _291_ = _018_;
    endcase
  assign \Mem[25]  = _291_;
  reg [15:0] _292_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _292_ = _088_;
      default:
        _292_ = _019_;
    endcase
  assign \Mem[26]  = _292_;
  reg [15:0] _293_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _293_ = _089_;
      default:
        _293_ = _020_;
    endcase
  assign \Mem[27]  = _293_;
  reg [15:0] _294_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _294_ = _090_;
      default:
        _294_ = _021_;
    endcase
  assign \Mem[28]  = _294_;
  reg [15:0] _295_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _295_ = _091_;
      default:
        _295_ = _022_;
    endcase
  assign \Mem[29]  = _295_;
  reg [15:0] _296_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _296_ = _092_;
      default:
        _296_ = _023_;
    endcase
  assign \Mem[2]  = _296_;
  reg [15:0] _297_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _297_ = _093_;
      default:
        _297_ = _024_;
    endcase
  assign \Mem[30]  = _297_;
  reg [15:0] _298_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _298_ = _094_;
      default:
        _298_ = _025_;
    endcase
  assign \Mem[31]  = _298_;
  reg [15:0] _299_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _299_ = _095_;
      default:
        _299_ = _026_;
    endcase
  assign \Mem[32]  = _299_;
  reg [15:0] _300_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _300_ = _096_;
      default:
        _300_ = _027_;
    endcase
  assign \Mem[33]  = _300_;
  reg [15:0] _301_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _301_ = _097_;
      default:
        _301_ = _028_;
    endcase
  assign \Mem[34]  = _301_;
  reg [15:0] _302_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _302_ = _098_;
      default:
        _302_ = _029_;
    endcase
  assign \Mem[35]  = _302_;
  reg [15:0] _303_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _303_ = _099_;
      default:
        _303_ = _030_;
    endcase
  assign \Mem[36]  = _303_;
  reg [15:0] _304_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _304_ = _100_;
      default:
        _304_ = _031_;
    endcase
  assign \Mem[37]  = _304_;
  reg [15:0] _305_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _305_ = _101_;
      default:
        _305_ = _032_;
    endcase
  assign \Mem[38]  = _305_;
  reg [15:0] _306_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _306_ = _102_;
      default:
        _306_ = _033_;
    endcase
  assign \Mem[39]  = _306_;
  reg [15:0] _307_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _307_ = _103_;
      default:
        _307_ = _034_;
    endcase
  assign \Mem[3]  = _307_;
  reg [15:0] _308_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _308_ = _104_;
      default:
        _308_ = _035_;
    endcase
  assign \Mem[40]  = _308_;
  reg [15:0] _309_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _309_ = _105_;
      default:
        _309_ = _036_;
    endcase
  assign \Mem[41]  = _309_;
  reg [15:0] _310_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _310_ = _106_;
      default:
        _310_ = _037_;
    endcase
  assign \Mem[42]  = _310_;
  reg [15:0] _311_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _311_ = _107_;
      default:
        _311_ = _038_;
    endcase
  assign \Mem[43]  = _311_;
  reg [15:0] _312_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _312_ = _108_;
      default:
        _312_ = _039_;
    endcase
  assign \Mem[44]  = _312_;
  reg [15:0] _313_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _313_ = _109_;
      default:
        _313_ = _040_;
    endcase
  assign \Mem[45]  = _313_;
  reg [15:0] _314_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _314_ = _110_;
      default:
        _314_ = _041_;
    endcase
  assign \Mem[46]  = _314_;
  reg [15:0] _315_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _315_ = _111_;
      default:
        _315_ = _042_;
    endcase
  assign \Mem[47]  = _315_;
  reg [15:0] _316_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _316_ = _112_;
      default:
        _316_ = _043_;
    endcase
  assign \Mem[48]  = _316_;
  reg [15:0] _317_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _317_ = _113_;
      default:
        _317_ = _044_;
    endcase
  assign \Mem[49]  = _317_;
  reg [15:0] _318_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _318_ = _114_;
      default:
        _318_ = _045_;
    endcase
  assign \Mem[4]  = _318_;
  reg [15:0] _319_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _319_ = _115_;
      default:
        _319_ = _046_;
    endcase
  assign \Mem[50]  = _319_;
  reg [15:0] _320_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _320_ = _116_;
      default:
        _320_ = _047_;
    endcase
  assign \Mem[51]  = _320_;
  reg [15:0] _321_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _321_ = _117_;
      default:
        _321_ = _048_;
    endcase
  assign \Mem[52]  = _321_;
  reg [15:0] _322_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _322_ = _118_;
      default:
        _322_ = _049_;
    endcase
  assign \Mem[53]  = _322_;
  reg [15:0] _323_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _323_ = _119_;
      default:
        _323_ = _050_;
    endcase
  assign \Mem[54]  = _323_;
  reg [15:0] _324_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _324_ = _120_;
      default:
        _324_ = _051_;
    endcase
  assign \Mem[55]  = _324_;
  reg [15:0] _325_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _325_ = _121_;
      default:
        _325_ = _052_;
    endcase
  assign \Mem[56]  = _325_;
  reg [15:0] _326_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _326_ = _122_;
      default:
        _326_ = _053_;
    endcase
  assign \Mem[57]  = _326_;
  reg [15:0] _327_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _327_ = _123_;
      default:
        _327_ = _054_;
    endcase
  assign \Mem[58]  = _327_;
  reg [15:0] _328_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _328_ = _124_;
      default:
        _328_ = _055_;
    endcase
  assign \Mem[59]  = _328_;
  reg [15:0] _329_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _329_ = _125_;
      default:
        _329_ = _056_;
    endcase
  assign \Mem[5]  = _329_;
  reg [15:0] _330_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _330_ = _126_;
      default:
        _330_ = _057_;
    endcase
  assign \Mem[60]  = _330_;
  reg [15:0] _331_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _331_ = _127_;
      default:
        _331_ = _058_;
    endcase
  assign \Mem[61]  = _331_;
  reg [15:0] _332_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _332_ = _128_;
      default:
        _332_ = _059_;
    endcase
  assign \Mem[62]  = _332_;
  reg [15:0] _333_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _333_ = _129_;
      default:
        _333_ = _060_;
    endcase
  assign _069_ = _333_;
  reg [15:0] _334_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _334_ = _130_;
      default:
        _334_ = _061_;
    endcase
  assign \Mem[6]  = _334_;
  reg [15:0] _335_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _335_ = _131_;
      default:
        _335_ = _062_;
    endcase
  assign \Mem[7]  = _335_;
  reg [15:0] _336_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _336_ = _132_;
      default:
        _336_ = _063_;
    endcase
  assign \Mem[8]  = _336_;
  reg [15:0] _337_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _337_ = _133_;
      default:
        _337_ = _064_;
    endcase
  assign \Mem[9]  = _337_;
  reg [0:0] _338_;
  (* parallel_case *)
  always @*
    casez (_136_)
      1'b1:
        _338_ = _068_;
      default:
        _338_ = _065_;
    endcase
  assign bug_a = _338_;
  reg [15:0] _339_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _339_ = 16'b0000000000000000;
      default:
        _339_ = _001_;
    endcase
  assign _070_ = _339_;
  reg [15:0] _340_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _340_ = 16'b0000000000000000;
      default:
        _340_ = _002_;
    endcase
  assign _071_ = _340_;
  reg [15:0] _341_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _341_ = 16'b0000000000000000;
      default:
        _341_ = _003_;
    endcase
  assign _072_ = _341_;
  reg [15:0] _342_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _342_ = 16'b0000000000000000;
      default:
        _342_ = _004_;
    endcase
  assign _073_ = _342_;
  reg [15:0] _343_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _343_ = 16'b0000000000000000;
      default:
        _343_ = _005_;
    endcase
  assign _074_ = _343_;
  reg [15:0] _344_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _344_ = 16'b0000000000000000;
      default:
        _344_ = _006_;
    endcase
  assign _075_ = _344_;
  reg [15:0] _345_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _345_ = 16'b0000000000000000;
      default:
        _345_ = _007_;
    endcase
  assign _076_ = _345_;
  reg [15:0] _346_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _346_ = 16'b0000000000000000;
      default:
        _346_ = _008_;
    endcase
  assign _077_ = _346_;
  reg [15:0] _347_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _347_ = 16'b0000000000000000;
      default:
        _347_ = _009_;
    endcase
  assign _078_ = _347_;
  reg [15:0] _348_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _348_ = 16'b0000000000000000;
      default:
        _348_ = _010_;
    endcase
  assign _079_ = _348_;
  reg [15:0] _349_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _349_ = 16'b0000000000000000;
      default:
        _349_ = _011_;
    endcase
  assign _080_ = _349_;
  reg [15:0] _350_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _350_ = 16'b0000000000000000;
      default:
        _350_ = _012_;
    endcase
  assign _081_ = _350_;
  reg [15:0] _351_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _351_ = 16'b0000000000000000;
      default:
        _351_ = _013_;
    endcase
  assign _082_ = _351_;
  reg [15:0] _352_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _352_ = 16'b0000000000000000;
      default:
        _352_ = _014_;
    endcase
  assign _083_ = _352_;
  reg [15:0] _353_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _353_ = 16'b0000000000000000;
      default:
        _353_ = _015_;
    endcase
  assign _084_ = _353_;
  reg [15:0] _354_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _354_ = 16'b0000000000000000;
      default:
        _354_ = _016_;
    endcase
  assign _085_ = _354_;
  reg [15:0] _355_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _355_ = 16'b0000000000000000;
      default:
        _355_ = _017_;
    endcase
  assign _086_ = _355_;
  reg [15:0] _356_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _356_ = 16'b0000000000000000;
      default:
        _356_ = _018_;
    endcase
  assign _087_ = _356_;
  reg [15:0] _357_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _357_ = 16'b0000000000000000;
      default:
        _357_ = _019_;
    endcase
  assign _088_ = _357_;
  reg [15:0] _358_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _358_ = 16'b0000000000000000;
      default:
        _358_ = _020_;
    endcase
  assign _089_ = _358_;
  reg [15:0] _359_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _359_ = 16'b0000000000000000;
      default:
        _359_ = _021_;
    endcase
  assign _090_ = _359_;
  reg [15:0] _360_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _360_ = 16'b0000000000000000;
      default:
        _360_ = _022_;
    endcase
  assign _091_ = _360_;
  reg [15:0] _361_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _361_ = 16'b0000000000000000;
      default:
        _361_ = _023_;
    endcase
  assign _092_ = _361_;
  reg [15:0] _362_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _362_ = 16'b0000000000000000;
      default:
        _362_ = _024_;
    endcase
  assign _093_ = _362_;
  reg [15:0] _363_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _363_ = 16'b0000000000000000;
      default:
        _363_ = _025_;
    endcase
  assign _094_ = _363_;
  reg [15:0] _364_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _364_ = 16'b0000000000000000;
      default:
        _364_ = _026_;
    endcase
  assign _095_ = _364_;
  reg [15:0] _365_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _365_ = 16'b0000000000000000;
      default:
        _365_ = _027_;
    endcase
  assign _096_ = _365_;
  reg [15:0] _366_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _366_ = 16'b0000000000000000;
      default:
        _366_ = _028_;
    endcase
  assign _097_ = _366_;
  reg [15:0] _367_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _367_ = 16'b0000000000000000;
      default:
        _367_ = _029_;
    endcase
  assign _098_ = _367_;
  reg [15:0] _368_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _368_ = 16'b0000000000000000;
      default:
        _368_ = _030_;
    endcase
  assign _099_ = _368_;
  reg [15:0] _369_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _369_ = 16'b0000000000000000;
      default:
        _369_ = _031_;
    endcase
  assign _100_ = _369_;
  reg [15:0] _370_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _370_ = 16'b0000000000000000;
      default:
        _370_ = _032_;
    endcase
  assign _101_ = _370_;
  reg [15:0] _371_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _371_ = 16'b0000000000000000;
      default:
        _371_ = _033_;
    endcase
  assign _102_ = _371_;
  reg [15:0] _372_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _372_ = 16'b0000000000000000;
      default:
        _372_ = _034_;
    endcase
  assign _103_ = _372_;
  reg [15:0] _373_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _373_ = 16'b0000000000000000;
      default:
        _373_ = _035_;
    endcase
  assign _104_ = _373_;
  reg [15:0] _374_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _374_ = 16'b0000000000000000;
      default:
        _374_ = _036_;
    endcase
  assign _105_ = _374_;
  reg [15:0] _375_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _375_ = 16'b0000000000000000;
      default:
        _375_ = _037_;
    endcase
  assign _106_ = _375_;
  reg [15:0] _376_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _376_ = 16'b0000000000000000;
      default:
        _376_ = _038_;
    endcase
  assign _107_ = _376_;
  reg [15:0] _377_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _377_ = 16'b0000000000000000;
      default:
        _377_ = _039_;
    endcase
  assign _108_ = _377_;
  reg [15:0] _378_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _378_ = 16'b0000000000000000;
      default:
        _378_ = _040_;
    endcase
  assign _109_ = _378_;
  reg [15:0] _379_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _379_ = 16'b0000000000000000;
      default:
        _379_ = _041_;
    endcase
  assign _110_ = _379_;
  reg [15:0] _380_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _380_ = 16'b0000000000000000;
      default:
        _380_ = _042_;
    endcase
  assign _111_ = _380_;
  reg [15:0] _381_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _381_ = 16'b0000000000000000;
      default:
        _381_ = _043_;
    endcase
  assign _112_ = _381_;
  reg [15:0] _382_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _382_ = 16'b0000000000000000;
      default:
        _382_ = _044_;
    endcase
  assign _113_ = _382_;
  reg [15:0] _383_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _383_ = 16'b0000000000000000;
      default:
        _383_ = _045_;
    endcase
  assign _114_ = _383_;
  reg [15:0] _384_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _384_ = 16'b0000000000000000;
      default:
        _384_ = _046_;
    endcase
  assign _115_ = _384_;
  reg [15:0] _385_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _385_ = 16'b0000000000000000;
      default:
        _385_ = _047_;
    endcase
  assign _116_ = _385_;
  reg [15:0] _386_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _386_ = 16'b0000000000000000;
      default:
        _386_ = _048_;
    endcase
  assign _117_ = _386_;
  reg [15:0] _387_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _387_ = 16'b0000000000000000;
      default:
        _387_ = _049_;
    endcase
  assign _118_ = _387_;
  reg [15:0] _388_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _388_ = 16'b0000000000000000;
      default:
        _388_ = _050_;
    endcase
  assign _119_ = _388_;
  reg [15:0] _389_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _389_ = 16'b0000000000000000;
      default:
        _389_ = _051_;
    endcase
  assign _120_ = _389_;
  reg [15:0] _390_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _390_ = 16'b0000000000000000;
      default:
        _390_ = _052_;
    endcase
  assign _121_ = _390_;
  reg [15:0] _391_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _391_ = 16'b0000000000000000;
      default:
        _391_ = _053_;
    endcase
  assign _122_ = _391_;
  reg [15:0] _392_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _392_ = 16'b0000000000000000;
      default:
        _392_ = _054_;
    endcase
  assign _123_ = _392_;
  reg [15:0] _393_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _393_ = 16'b0000000000000000;
      default:
        _393_ = _055_;
    endcase
  assign _124_ = _393_;
  reg [15:0] _394_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _394_ = 16'b0000000000000000;
      default:
        _394_ = _056_;
    endcase
  assign _125_ = _394_;
  reg [15:0] _395_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _395_ = 16'b0000000000000000;
      default:
        _395_ = _057_;
    endcase
  assign _126_ = _395_;
  reg [15:0] _396_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _396_ = 16'b0000000000000000;
      default:
        _396_ = _058_;
    endcase
  assign _127_ = _396_;
  reg [15:0] _397_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _397_ = 16'b0000000000000000;
      default:
        _397_ = _059_;
    endcase
  assign _128_ = _397_;
  reg [15:0] _398_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _398_ = 16'b0000000000000000;
      default:
        _398_ = _060_;
    endcase
  assign _129_ = _398_;
  reg [15:0] _399_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _399_ = 16'b0000000000000000;
      default:
        _399_ = _061_;
    endcase
  assign _130_ = _399_;
  reg [15:0] _400_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _400_ = 16'b0000000000000000;
      default:
        _400_ = _062_;
    endcase
  assign _131_ = _400_;
  reg [15:0] _401_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _401_ = 16'b0000000000000000;
      default:
        _401_ = _063_;
    endcase
  assign _132_ = _401_;
  reg [15:0] _402_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _402_ = 16'b0000000000000000;
      default:
        _402_ = _064_;
    endcase
  assign _133_ = _402_;
  reg [0:0] _403_;
  (* parallel_case *)
  always @*
    casez (_065_)
      1'b1:
        _403_ = 1'b0;
      default:
        _403_ = _065_;
    endcase
  assign _068_ = _403_;
  reg [15:0] _404_;
  (* parallel_case *)
  always @*
    casez (WE)
      1'b1:
        _404_ = 16'b0000000000000000;
      default:
        _404_ = _069_;
    endcase
  assign \Mem[63]  = _404_;
  reg [15:0] _405_;
  (* parallel_case *)
  always @*
    casez ({ _158_, _157_, _156_, _155_, _154_, _153_, _152_, _151_, _150_, _149_, _148_, _147_, _146_, _145_, _144_, _143_, _142_, _141_, _177_, _176_, _175_, _174_, _173_, _172_, _171_, _170_, _169_, _168_, _167_, _166_, _165_, _164_, _163_, _162_, _161_, _160_, _159_, _178_, _179_, _180_, _181_, _182_, _183_, _184_, _185_, _186_, _187_, _188_, _189_, _190_, _191_, _192_, _193_, _194_, _195_, _196_, _197_, _198_, _199_, _200_, _201_, _202_, _203_ })
      63'b??????????????????????????????????????????????????????????????1:
        _405_ = \Mem[62] ;
      63'b?????????????????????????????????????????????????????????????1?:
        _405_ = \Mem[61] ;
      63'b????????????????????????????????????????????????????????????1??:
        _405_ = \Mem[60] ;
      63'b???????????????????????????????????????????????????????????1???:
        _405_ = \Mem[59] ;
      63'b??????????????????????????????????????????????????????????1????:
        _405_ = \Mem[58] ;
      63'b?????????????????????????????????????????????????????????1?????:
        _405_ = \Mem[57] ;
      63'b????????????????????????????????????????????????????????1??????:
        _405_ = \Mem[56] ;
      63'b???????????????????????????????????????????????????????1???????:
        _405_ = \Mem[55] ;
      63'b??????????????????????????????????????????????????????1????????:
        _405_ = \Mem[54] ;
      63'b?????????????????????????????????????????????????????1?????????:
        _405_ = \Mem[53] ;
      63'b????????????????????????????????????????????????????1??????????:
        _405_ = \Mem[52] ;
      63'b???????????????????????????????????????????????????1???????????:
        _405_ = \Mem[51] ;
      63'b??????????????????????????????????????????????????1????????????:
        _405_ = \Mem[50] ;
      63'b?????????????????????????????????????????????????1?????????????:
        _405_ = \Mem[49] ;
      63'b????????????????????????????????????????????????1??????????????:
        _405_ = \Mem[48] ;
      63'b???????????????????????????????????????????????1???????????????:
        _405_ = \Mem[47] ;
      63'b??????????????????????????????????????????????1????????????????:
        _405_ = \Mem[46] ;
      63'b?????????????????????????????????????????????1?????????????????:
        _405_ = \Mem[45] ;
      63'b????????????????????????????????????????????1??????????????????:
        _405_ = \Mem[44] ;
      63'b???????????????????????????????????????????1???????????????????:
        _405_ = \Mem[43] ;
      63'b??????????????????????????????????????????1????????????????????:
        _405_ = \Mem[42] ;
      63'b?????????????????????????????????????????1?????????????????????:
        _405_ = \Mem[41] ;
      63'b????????????????????????????????????????1??????????????????????:
        _405_ = \Mem[40] ;
      63'b???????????????????????????????????????1???????????????????????:
        _405_ = \Mem[39] ;
      63'b??????????????????????????????????????1????????????????????????:
        _405_ = \Mem[38] ;
      63'b?????????????????????????????????????1?????????????????????????:
        _405_ = \Mem[37] ;
      63'b????????????????????????????????????1??????????????????????????:
        _405_ = \Mem[36] ;
      63'b???????????????????????????????????1???????????????????????????:
        _405_ = \Mem[35] ;
      63'b??????????????????????????????????1????????????????????????????:
        _405_ = \Mem[34] ;
      63'b?????????????????????????????????1?????????????????????????????:
        _405_ = \Mem[33] ;
      63'b????????????????????????????????1??????????????????????????????:
        _405_ = \Mem[32] ;
      63'b???????????????????????????????1???????????????????????????????:
        _405_ = \Mem[31] ;
      63'b??????????????????????????????1????????????????????????????????:
        _405_ = \Mem[30] ;
      63'b?????????????????????????????1?????????????????????????????????:
        _405_ = \Mem[29] ;
      63'b????????????????????????????1??????????????????????????????????:
        _405_ = \Mem[28] ;
      63'b???????????????????????????1???????????????????????????????????:
        _405_ = \Mem[27] ;
      63'b??????????????????????????1????????????????????????????????????:
        _405_ = \Mem[26] ;
      63'b?????????????????????????1?????????????????????????????????????:
        _405_ = \Mem[25] ;
      63'b????????????????????????1??????????????????????????????????????:
        _405_ = \Mem[24] ;
      63'b???????????????????????1???????????????????????????????????????:
        _405_ = \Mem[23] ;
      63'b??????????????????????1????????????????????????????????????????:
        _405_ = \Mem[22] ;
      63'b?????????????????????1?????????????????????????????????????????:
        _405_ = \Mem[21] ;
      63'b????????????????????1??????????????????????????????????????????:
        _405_ = \Mem[20] ;
      63'b???????????????????1???????????????????????????????????????????:
        _405_ = \Mem[19] ;
      63'b??????????????????1????????????????????????????????????????????:
        _405_ = \Mem[18] ;
      63'b?????????????????1?????????????????????????????????????????????:
        _405_ = \Mem[17] ;
      63'b????????????????1??????????????????????????????????????????????:
        _405_ = \Mem[16] ;
      63'b???????????????1???????????????????????????????????????????????:
        _405_ = \Mem[15] ;
      63'b??????????????1????????????????????????????????????????????????:
        _405_ = \Mem[14] ;
      63'b?????????????1?????????????????????????????????????????????????:
        _405_ = \Mem[13] ;
      63'b????????????1??????????????????????????????????????????????????:
        _405_ = \Mem[12] ;
      63'b???????????1???????????????????????????????????????????????????:
        _405_ = \Mem[11] ;
      63'b??????????1????????????????????????????????????????????????????:
        _405_ = \Mem[10] ;
      63'b?????????1?????????????????????????????????????????????????????:
        _405_ = \Mem[9] ;
      63'b????????1??????????????????????????????????????????????????????:
        _405_ = \Mem[8] ;
      63'b???????1???????????????????????????????????????????????????????:
        _405_ = \Mem[7] ;
      63'b??????1????????????????????????????????????????????????????????:
        _405_ = \Mem[6] ;
      63'b?????1?????????????????????????????????????????????????????????:
        _405_ = \Mem[5] ;
      63'b????1??????????????????????????????????????????????????????????:
        _405_ = \Mem[4] ;
      63'b???1???????????????????????????????????????????????????????????:
        _405_ = \Mem[3] ;
      63'b??1????????????????????????????????????????????????????????????:
        _405_ = \Mem[2] ;
      63'b?1?????????????????????????????????????????????????????????????:
        _405_ = \Mem[1] ;
      63'b1??????????????????????????????????????????????????????????????:
        _405_ = \Mem[0] ;
      default:
        _405_ = \Mem[63] ;
    endcase
  assign _000_ = _405_;
  reg [15:0] _406_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _406_ = _067_;
      default:
        _406_ = \Mem[0] ;
    endcase
  assign _001_ = _406_;
  reg [15:0] _407_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _407_ = _067_;
      default:
        _407_ = \Mem[10] ;
    endcase
  assign _002_ = _407_;
  reg [15:0] _408_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _408_ = _067_;
      default:
        _408_ = \Mem[11] ;
    endcase
  assign _003_ = _408_;
  reg [15:0] _409_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _409_ = _067_;
      default:
        _409_ = \Mem[12] ;
    endcase
  assign _004_ = _409_;
  reg [15:0] _410_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _410_ = _067_;
      default:
        _410_ = \Mem[13] ;
    endcase
  assign _005_ = _410_;
  reg [15:0] _411_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _411_ = _067_;
      default:
        _411_ = \Mem[14] ;
    endcase
  assign _006_ = _411_;
  reg [15:0] _412_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _412_ = _067_;
      default:
        _412_ = \Mem[15] ;
    endcase
  assign _007_ = _412_;
  reg [15:0] _413_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _413_ = _067_;
      default:
        _413_ = \Mem[16] ;
    endcase
  assign _008_ = _413_;
  reg [15:0] _414_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _414_ = _067_;
      default:
        _414_ = \Mem[17] ;
    endcase
  assign _009_ = _414_;
  reg [15:0] _415_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _415_ = _067_;
      default:
        _415_ = \Mem[18] ;
    endcase
  assign _010_ = _415_;
  reg [15:0] _416_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _416_ = _067_;
      default:
        _416_ = \Mem[19] ;
    endcase
  assign _011_ = _416_;
  reg [15:0] _417_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _417_ = _067_;
      default:
        _417_ = \Mem[1] ;
    endcase
  assign _012_ = _417_;
  reg [15:0] _418_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _418_ = _067_;
      default:
        _418_ = \Mem[20] ;
    endcase
  assign _013_ = _418_;
  reg [15:0] _419_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _419_ = _067_;
      default:
        _419_ = \Mem[21] ;
    endcase
  assign _014_ = _419_;
  reg [15:0] _420_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _420_ = _067_;
      default:
        _420_ = \Mem[22] ;
    endcase
  assign _015_ = _420_;
  reg [15:0] _421_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _421_ = _067_;
      default:
        _421_ = \Mem[23] ;
    endcase
  assign _016_ = _421_;
  reg [15:0] _422_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _422_ = _067_;
      default:
        _422_ = \Mem[24] ;
    endcase
  assign _017_ = _422_;
  reg [15:0] _423_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _423_ = _067_;
      default:
        _423_ = \Mem[25] ;
    endcase
  assign _018_ = _423_;
  reg [15:0] _424_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _424_ = _067_;
      default:
        _424_ = \Mem[26] ;
    endcase
  assign _019_ = _424_;
  reg [15:0] _425_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _425_ = _067_;
      default:
        _425_ = \Mem[27] ;
    endcase
  assign _020_ = _425_;
  reg [15:0] _426_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _426_ = _067_;
      default:
        _426_ = \Mem[28] ;
    endcase
  assign _021_ = _426_;
  reg [15:0] _427_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _427_ = _067_;
      default:
        _427_ = \Mem[29] ;
    endcase
  assign _022_ = _427_;
  reg [15:0] _428_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _428_ = _067_;
      default:
        _428_ = \Mem[2] ;
    endcase
  assign _023_ = _428_;
  reg [15:0] _429_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _429_ = _067_;
      default:
        _429_ = \Mem[30] ;
    endcase
  assign _024_ = _429_;
  reg [15:0] _430_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _430_ = _067_;
      default:
        _430_ = \Mem[31] ;
    endcase
  assign _025_ = _430_;
  reg [15:0] _431_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _431_ = _067_;
      default:
        _431_ = \Mem[32] ;
    endcase
  assign _026_ = _431_;
  reg [15:0] _432_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _432_ = _067_;
      default:
        _432_ = \Mem[33] ;
    endcase
  assign _027_ = _432_;
  reg [15:0] _433_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _433_ = _067_;
      default:
        _433_ = \Mem[34] ;
    endcase
  assign _028_ = _433_;
  reg [15:0] _434_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _434_ = _067_;
      default:
        _434_ = \Mem[35] ;
    endcase
  assign _029_ = _434_;
  reg [15:0] _435_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _435_ = _067_;
      default:
        _435_ = \Mem[36] ;
    endcase
  assign _030_ = _435_;
  reg [15:0] _436_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _436_ = _067_;
      default:
        _436_ = \Mem[37] ;
    endcase
  assign _031_ = _436_;
  reg [15:0] _437_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _437_ = _067_;
      default:
        _437_ = \Mem[38] ;
    endcase
  assign _032_ = _437_;
  reg [15:0] _438_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _438_ = _067_;
      default:
        _438_ = \Mem[39] ;
    endcase
  assign _033_ = _438_;
  reg [15:0] _439_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _439_ = _067_;
      default:
        _439_ = \Mem[3] ;
    endcase
  assign _034_ = _439_;
  reg [15:0] _440_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _440_ = _067_;
      default:
        _440_ = \Mem[40] ;
    endcase
  assign _035_ = _440_;
  reg [15:0] _441_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _441_ = _067_;
      default:
        _441_ = \Mem[41] ;
    endcase
  assign _036_ = _441_;
  reg [15:0] _442_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _442_ = _067_;
      default:
        _442_ = \Mem[42] ;
    endcase
  assign _037_ = _442_;
  reg [15:0] _443_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _443_ = _067_;
      default:
        _443_ = \Mem[43] ;
    endcase
  assign _038_ = _443_;
  reg [15:0] _444_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _444_ = _067_;
      default:
        _444_ = \Mem[44] ;
    endcase
  assign _039_ = _444_;
  reg [15:0] _445_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _445_ = _067_;
      default:
        _445_ = \Mem[45] ;
    endcase
  assign _040_ = _445_;
  reg [15:0] _446_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _446_ = _067_;
      default:
        _446_ = \Mem[46] ;
    endcase
  assign _041_ = _446_;
  reg [15:0] _447_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _447_ = _067_;
      default:
        _447_ = \Mem[47] ;
    endcase
  assign _042_ = _447_;
  reg [15:0] _448_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _448_ = _067_;
      default:
        _448_ = \Mem[48] ;
    endcase
  assign _043_ = _448_;
  reg [15:0] _449_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _449_ = _067_;
      default:
        _449_ = \Mem[49] ;
    endcase
  assign _044_ = _449_;
  reg [15:0] _450_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _450_ = _067_;
      default:
        _450_ = \Mem[4] ;
    endcase
  assign _045_ = _450_;
  reg [15:0] _451_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _451_ = _067_;
      default:
        _451_ = \Mem[50] ;
    endcase
  assign _046_ = _451_;
  reg [15:0] _452_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _452_ = _067_;
      default:
        _452_ = \Mem[51] ;
    endcase
  assign _047_ = _452_;
  reg [15:0] _453_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _453_ = _067_;
      default:
        _453_ = \Mem[52] ;
    endcase
  assign _048_ = _453_;
  reg [15:0] _454_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _454_ = _067_;
      default:
        _454_ = \Mem[53] ;
    endcase
  assign _049_ = _454_;
  reg [15:0] _455_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _455_ = _067_;
      default:
        _455_ = \Mem[54] ;
    endcase
  assign _050_ = _455_;
  reg [15:0] _456_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _456_ = _067_;
      default:
        _456_ = \Mem[55] ;
    endcase
  assign _051_ = _456_;
  reg [15:0] _457_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _457_ = _067_;
      default:
        _457_ = \Mem[56] ;
    endcase
  assign _052_ = _457_;
  reg [15:0] _458_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _458_ = _067_;
      default:
        _458_ = \Mem[57] ;
    endcase
  assign _053_ = _458_;
  reg [15:0] _459_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _459_ = _067_;
      default:
        _459_ = \Mem[58] ;
    endcase
  assign _054_ = _459_;
  reg [15:0] _460_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _460_ = _067_;
      default:
        _460_ = \Mem[59] ;
    endcase
  assign _055_ = _460_;
  reg [15:0] _461_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _461_ = _067_;
      default:
        _461_ = \Mem[5] ;
    endcase
  assign _056_ = _461_;
  reg [15:0] _462_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _462_ = _067_;
      default:
        _462_ = \Mem[60] ;
    endcase
  assign _057_ = _462_;
  reg [15:0] _463_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _463_ = _067_;
      default:
        _463_ = \Mem[61] ;
    endcase
  assign _058_ = _463_;
  reg [15:0] _464_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _464_ = _067_;
      default:
        _464_ = \Mem[62] ;
    endcase
  assign _059_ = _464_;
  reg [15:0] _465_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _465_ = _067_;
      default:
        _465_ = \Mem[63] ;
    endcase
  assign _060_ = _465_;
  reg [15:0] _466_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _466_ = _067_;
      default:
        _466_ = \Mem[6] ;
    endcase
  assign _061_ = _466_;
  reg [15:0] _467_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _467_ = _067_;
      default:
        _467_ = \Mem[7] ;
    endcase
  assign _062_ = _467_;
  reg [15:0] _468_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _468_ = _067_;
      default:
        _468_ = \Mem[8] ;
    endcase
  assign _063_ = _468_;
  reg [15:0] _469_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _469_ = _067_;
      default:
        _469_ = \Mem[9] ;
    endcase
  assign _064_ = _469_;
  reg [0:0] _470_;
  (* parallel_case *)
  always @*
    casez (_134_)
      1'b1:
        _470_ = _066_;
      default:
        _470_ = bug_a;
    endcase
  assign _065_ = _470_;
  reg [15:0] _471_;
  (* parallel_case *)
  always @*
    casez (_135_)
      1'b1:
        _471_ = 16'b0000000000000000;
      default:
        _471_ = Data;
    endcase
  assign _067_ = _471_;
  reg [0:0] _472_;
  (* parallel_case *)
  always @*
    casez (_135_)
      1'b1:
        _472_ = 1'b1;
      default:
        _472_ = bug_a;
    endcase
  assign _066_ = _472_;
  reg [15:0] _473_;
  (* src = "design.sv:14" *)
  (* parallel_case *)
  always @*
    casez (OE)
      1'b1:
        _473_ = 16'bzzzzzzzzzzzzzzzz;
      default:
        _473_ = _000_;
    endcase
  assign Data = _473_;
endmodule
